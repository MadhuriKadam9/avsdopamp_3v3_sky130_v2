* SPICE3 file created from res.ext - technology: sky130A

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 b a SUB sky130_fd_pr__res_generic_nd w=20 l=50

Va a 0 dc 3.3

Vb b 0 dc 0

.tran 0.1us 20us
.control
run

plot V(a)/(-Va#branch)

.endc

.end
