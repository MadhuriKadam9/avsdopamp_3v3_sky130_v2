magic
tech sky130A
timestamp 1628848859
<< nwell >>
rect -634 183 7076 1735
rect -634 -1455 7076 -196
<< nmos >>
rect 1505 -2003 2504 -1947
rect 3208 -2010 4207 -1954
<< pmos >>
rect 2380 652 3384 700
rect 80 -555 2592 -503
rect 3212 -547 5724 -495
<< ndiff >>
rect 1505 -1812 2504 -1746
rect 1505 -1887 1569 -1812
rect 1793 -1887 2208 -1812
rect 2432 -1887 2504 -1812
rect 1505 -1947 2504 -1887
rect 3208 -1819 4207 -1753
rect 3208 -1894 3272 -1819
rect 3496 -1894 3911 -1819
rect 4135 -1894 4207 -1819
rect 3208 -1954 4207 -1894
rect 1505 -2078 2504 -2003
rect 1505 -2171 1573 -2078
rect 1797 -2171 2189 -2078
rect 2413 -2171 2504 -2078
rect 1505 -2201 2504 -2171
rect 3208 -2085 4207 -2010
rect 3208 -2178 3276 -2085
rect 3500 -2178 3892 -2085
rect 4116 -2178 4207 -2085
rect 3208 -2208 4207 -2178
<< pdiff >>
rect 2380 996 3384 1058
rect 2380 808 2432 996
rect 2632 984 3384 996
rect 2632 808 3152 984
rect 2380 796 3152 808
rect 3352 796 3384 984
rect 2380 700 3384 796
rect 2380 580 3384 652
rect 2380 568 3144 580
rect 2380 380 2432 568
rect 2632 392 3144 568
rect 3344 392 3384 580
rect 2632 380 3384 392
rect 2380 341 3384 380
rect 80 -344 2592 -297
rect 80 -356 1004 -344
rect 80 -463 122 -356
rect 674 -451 1004 -356
rect 1556 -348 2592 -344
rect 1556 -451 1997 -348
rect 2549 -451 2592 -348
rect 674 -463 2592 -451
rect 80 -503 2592 -463
rect 3212 -336 5724 -289
rect 3212 -348 4136 -336
rect 3212 -455 3254 -348
rect 3806 -443 4136 -348
rect 4688 -340 5724 -336
rect 4688 -443 5129 -340
rect 5681 -443 5724 -340
rect 3806 -455 5724 -443
rect 3212 -495 5724 -455
rect 80 -610 2592 -555
rect 80 -614 2001 -610
rect 80 -717 122 -614
rect 674 -618 2001 -614
rect 674 -717 1012 -618
rect 80 -725 1012 -717
rect 1564 -713 2001 -618
rect 2553 -713 2592 -610
rect 1564 -725 2592 -713
rect 80 -757 2592 -725
rect 3212 -602 5724 -547
rect 3212 -606 5133 -602
rect 3212 -709 3254 -606
rect 3806 -610 5133 -606
rect 3806 -709 4144 -610
rect 3212 -717 4144 -709
rect 4696 -705 5133 -610
rect 5685 -705 5724 -602
rect 4696 -717 5724 -705
rect 3212 -749 5724 -717
<< ndiffc >>
rect 1569 -1887 1793 -1812
rect 2208 -1887 2432 -1812
rect 3272 -1894 3496 -1819
rect 3911 -1894 4135 -1819
rect 1573 -2171 1797 -2078
rect 2189 -2171 2413 -2078
rect 3276 -2178 3500 -2085
rect 3892 -2178 4116 -2085
<< pdiffc >>
rect 2432 808 2632 996
rect 3152 796 3352 984
rect 2432 380 2632 568
rect 3144 392 3344 580
rect 122 -463 674 -356
rect 1004 -451 1556 -344
rect 1997 -451 2549 -348
rect 3254 -455 3806 -348
rect 4136 -443 4688 -336
rect 5129 -443 5681 -340
rect 122 -717 674 -614
rect 1012 -725 1564 -618
rect 2001 -713 2553 -610
rect 3254 -709 3806 -606
rect 4144 -717 4696 -610
rect 5133 -705 5685 -602
<< psubdiff >>
rect 1498 -2276 2500 -2249
rect 1498 -2392 1561 -2276
rect 1789 -2279 2500 -2276
rect 1789 -2392 2189 -2279
rect 1498 -2395 2189 -2392
rect 2417 -2395 2500 -2279
rect 1498 -2451 2500 -2395
rect 3201 -2283 4203 -2256
rect 3201 -2399 3264 -2283
rect 3492 -2286 4203 -2283
rect 3492 -2399 3892 -2286
rect 3201 -2402 3892 -2399
rect 4120 -2402 4203 -2286
rect 3201 -2452 4203 -2402
<< nsubdiff >>
rect 2380 1387 3384 1441
rect 2380 1383 3116 1387
rect 2380 1195 2444 1383
rect 2644 1199 3116 1383
rect 3316 1199 3384 1387
rect 2644 1195 3384 1199
rect 2380 1098 3384 1195
<< psubdiffcont >>
rect 1561 -2392 1789 -2276
rect 2189 -2395 2417 -2279
rect 3264 -2399 3492 -2283
rect 3892 -2402 4120 -2286
<< nsubdiffcont >>
rect 2444 1195 2644 1383
rect 3116 1199 3316 1387
<< poly >>
rect 2119 688 2380 700
rect 2119 596 2156 688
rect 2256 652 2380 688
rect 3384 652 3475 700
rect 2256 596 2296 652
rect 2119 559 2296 596
rect -313 -424 -66 -392
rect -313 -575 -281 -424
rect -90 -471 -66 -424
rect -90 -503 29 -471
rect 5886 -392 6133 -384
rect 5886 -455 5934 -392
rect 5782 -495 5934 -455
rect -90 -555 80 -503
rect 2592 -555 2635 -503
rect 3161 -547 3212 -495
rect 5724 -543 5934 -495
rect 6125 -543 6133 -392
rect 5724 -547 6133 -543
rect -90 -575 29 -555
rect -313 -591 29 -575
rect -313 -647 -66 -591
rect 5782 -575 6133 -547
rect 5886 -639 6133 -575
rect 2554 -1933 3148 -1910
rect 2554 -1947 2719 -1933
rect 1397 -2003 1505 -1947
rect 2504 -1982 2719 -1947
rect 2768 -1954 3148 -1933
rect 2768 -1982 3208 -1954
rect 2504 -2001 3208 -1982
rect 2504 -2003 2601 -2001
rect 3100 -2010 3208 -2001
rect 4207 -2010 4304 -1954
<< polycont >>
rect 2156 596 2256 688
rect -281 -575 -90 -424
rect 5934 -543 6125 -392
rect 2719 -1982 2768 -1933
<< locali >>
rect 2381 1387 3387 1447
rect 2381 1383 3112 1387
rect 2381 1195 2444 1383
rect 2644 1203 3112 1383
rect 2644 1199 3116 1203
rect 3316 1199 3387 1387
rect 2644 1195 3387 1199
rect 2381 996 3387 1195
rect 2381 812 2428 996
rect 2632 984 3387 996
rect 2381 808 2432 812
rect 2632 808 3152 984
rect 3352 980 3387 984
rect 2381 796 3152 808
rect 3356 796 3387 980
rect 2381 728 3387 796
rect 2115 688 2292 696
rect 2115 596 2156 688
rect 2256 596 2292 688
rect 2115 555 2292 596
rect 2381 580 3383 620
rect 2381 568 3144 580
rect 2381 380 2432 568
rect 2632 392 3144 568
rect 3344 392 3383 580
rect 2632 380 3383 392
rect 2381 364 3383 380
rect 2365 332 3439 364
rect 2365 244 2592 332
rect 2323 -196 2592 244
rect 3212 252 3439 332
rect 3212 183 3487 252
rect 3218 -196 3487 183
rect 2300 -247 2592 -196
rect 2300 -292 2587 -247
rect 90 -336 2587 -292
rect 3216 -284 3503 -196
rect 3216 -336 5717 -284
rect 90 -344 2585 -336
rect 90 -356 1004 -344
rect -321 -424 -50 -392
rect -321 -575 -281 -424
rect -90 -575 -50 -424
rect 90 -463 122 -356
rect 674 -451 1004 -356
rect 1556 -348 2585 -344
rect 1556 -451 1997 -348
rect 2549 -451 2585 -348
rect 674 -463 2585 -451
rect 90 -483 2585 -463
rect 3222 -348 4136 -336
rect 3222 -455 3254 -348
rect 3806 -443 4136 -348
rect 4688 -340 5717 -336
rect 4688 -443 5129 -340
rect 5681 -443 5717 -340
rect 3806 -455 5717 -443
rect 3222 -475 5717 -455
rect 5870 -392 6141 -384
rect 5870 -543 5934 -392
rect 6125 -543 6141 -392
rect -321 -647 -50 -575
rect 94 -610 2589 -570
rect 94 -614 2001 -610
rect 94 -717 122 -614
rect 674 -618 2001 -614
rect 674 -717 1012 -618
rect 94 -725 1012 -717
rect 1564 -713 2001 -618
rect 2553 -713 2589 -610
rect 1564 -725 2589 -713
rect 94 -761 2589 -725
rect 3226 -602 5721 -562
rect 3226 -606 5133 -602
rect 3226 -709 3254 -606
rect 3806 -610 5133 -606
rect 3806 -709 4144 -610
rect 3226 -717 4144 -709
rect 4696 -705 5133 -610
rect 5685 -705 5721 -602
rect 5870 -639 6141 -543
rect 4696 -717 5721 -705
rect 3226 -753 5721 -717
rect 2340 -876 2499 -761
rect 2332 -989 2499 -876
rect 3296 -878 3440 -753
rect 3296 -934 3452 -878
rect 2332 -1523 2486 -989
rect 2332 -1595 2821 -1523
rect 2332 -1632 2828 -1595
rect 2332 -1779 2486 -1632
rect 1535 -1801 2486 -1779
rect 1535 -1812 2477 -1801
rect 1535 -1887 1569 -1812
rect 1793 -1887 2208 -1812
rect 2432 -1887 2477 -1812
rect 1535 -1913 2477 -1887
rect 2700 -1933 2828 -1632
rect 3298 -1786 3452 -934
rect 3238 -1819 4180 -1786
rect 3238 -1894 3272 -1819
rect 3496 -1894 3911 -1819
rect 4135 -1894 4180 -1819
rect 3238 -1920 4180 -1894
rect 2700 -1982 2719 -1933
rect 2768 -1982 2828 -1933
rect 2700 -2008 2828 -1982
rect 1524 -2078 2477 -2029
rect 1524 -2171 1573 -2078
rect 1797 -2171 2189 -2078
rect 2413 -2171 2477 -2078
rect 1524 -2276 2477 -2171
rect 1524 -2396 1561 -2276
rect 1789 -2279 2477 -2276
rect 1790 -2395 2189 -2279
rect 2417 -2395 2477 -2279
rect 1790 -2396 2193 -2395
rect 2411 -2396 2477 -2395
rect 1524 -2429 2477 -2396
rect 3227 -2085 4180 -2036
rect 3227 -2178 3276 -2085
rect 3500 -2178 3892 -2085
rect 4116 -2178 4180 -2085
rect 3227 -2283 4180 -2178
rect 3227 -2399 3264 -2283
rect 3492 -2286 4180 -2283
rect 3497 -2396 3889 -2286
rect 3492 -2399 3892 -2396
rect 3227 -2402 3892 -2399
rect 4120 -2402 4180 -2286
rect 3227 -2436 4180 -2402
<< viali >>
rect 2444 1195 2640 1383
rect 3112 1203 3116 1387
rect 3116 1203 3316 1387
rect 2428 812 2432 996
rect 2432 812 2632 996
rect 3152 796 3352 980
rect 3352 796 3356 980
rect 1561 -2392 1789 -2279
rect 1789 -2392 1790 -2279
rect 1561 -2396 1790 -2392
rect 2193 -2395 2411 -2279
rect 2193 -2396 2411 -2395
rect 3268 -2396 3492 -2286
rect 3492 -2396 3497 -2286
rect 3889 -2396 3892 -2286
rect 3892 -2396 4118 -2286
<< metal1 >>
rect 2341 1387 3415 1431
rect 2341 1383 3112 1387
rect 2341 1195 2444 1383
rect 2640 1203 3112 1383
rect 3316 1203 3415 1387
rect 2640 1195 3415 1203
rect 2341 996 3415 1195
rect 2341 812 2428 996
rect 2632 980 3415 996
rect 2632 812 3152 980
rect 2341 796 3152 812
rect 3356 796 3415 980
rect 2341 756 3415 796
rect 1444 -2049 2554 -2042
rect 1435 -2279 4258 -2049
rect 1435 -2396 1561 -2279
rect 1790 -2396 2193 -2279
rect 2411 -2286 4258 -2279
rect 2411 -2396 3268 -2286
rect 3497 -2396 3889 -2286
rect 4118 -2396 4258 -2286
rect 1435 -2420 4258 -2396
rect 1444 -2426 2554 -2420
rect 3148 -2433 4258 -2420
<< labels >>
rlabel locali 2787 -1993 2806 -1929 1 vg
rlabel metal1 1819 -2413 1875 -2275 1 gnd
rlabel locali 3354 -1615 3404 -1483 1 vo
rlabel locali -281 -647 -106 -591 1 vinp
rlabel locali 5941 -631 6116 -575 1 vinm
rlabel metal1 2459 1098 2636 1162 1 vdd
rlabel locali 2148 559 2256 588 1 vbias
<< end >>
