magic
tech sky130A
timestamp 1629199385
<< nwell >>
rect 6930 3789 9989 3797
rect -738 2237 9989 3789
rect 6930 2227 9989 2237
rect -738 1128 6196 1858
rect -738 599 3981 1128
<< nmos >>
rect 6948 1499 9468 1552
rect 1401 51 2400 107
rect 3104 44 4103 100
<< pmos >>
rect 2276 2706 3280 2754
rect 7848 2722 8864 2772
rect -24 1499 2488 1551
rect 3108 1507 5620 1559
<< ndiff >>
rect 6948 1729 9468 1757
rect 6948 1724 8920 1729
rect 6948 1626 7006 1724
rect 7481 1719 8920 1724
rect 7481 1626 7951 1719
rect 6948 1621 7951 1626
rect 8426 1631 8920 1719
rect 9395 1631 9468 1729
rect 8426 1621 9468 1631
rect 6948 1552 9468 1621
rect 6948 1421 9468 1499
rect 6948 1411 7946 1421
rect 6948 1313 7001 1411
rect 7476 1323 7946 1411
rect 8421 1323 8920 1421
rect 9395 1323 9468 1421
rect 7476 1313 9468 1323
rect 6948 1281 9468 1313
rect 1401 242 2400 308
rect 1401 167 1465 242
rect 1689 167 2104 242
rect 2328 167 2400 242
rect 1401 107 2400 167
rect 3104 235 4103 301
rect 3104 160 3168 235
rect 3392 160 3807 235
rect 4031 160 4103 235
rect 3104 100 4103 160
rect 1401 -24 2400 51
rect 1401 -117 1469 -24
rect 1693 -117 2085 -24
rect 2309 -117 2400 -24
rect 1401 -147 2400 -117
rect 3104 -31 4103 44
rect 3104 -124 3172 -31
rect 3396 -124 3788 -31
rect 4012 -124 4103 -31
rect 3104 -154 4103 -124
<< pdiff >>
rect 2276 3050 3280 3112
rect 2276 2862 2328 3050
rect 2528 3038 3280 3050
rect 2528 2862 3048 3038
rect 2276 2850 3048 2862
rect 3248 2850 3280 3038
rect 7848 3030 8864 3096
rect 2276 2754 3280 2850
rect 7848 2883 7910 3030
rect 8244 2883 8462 3030
rect 8796 2883 8864 3030
rect 7848 2772 8864 2883
rect 2276 2634 3280 2706
rect 2276 2622 3040 2634
rect 2276 2434 2328 2622
rect 2528 2446 3040 2622
rect 3240 2446 3280 2634
rect 2528 2434 3280 2446
rect 2276 2395 3280 2434
rect 7848 2625 8864 2722
rect 7848 2610 8477 2625
rect 7848 2463 7910 2610
rect 8244 2478 8477 2610
rect 8811 2478 8864 2625
rect 8244 2463 8864 2478
rect 7848 2405 8864 2463
rect -24 1710 2488 1757
rect -24 1698 900 1710
rect -24 1591 18 1698
rect 570 1603 900 1698
rect 1452 1706 2488 1710
rect 1452 1603 1893 1706
rect 2445 1603 2488 1706
rect 570 1591 2488 1603
rect -24 1551 2488 1591
rect 3108 1718 5620 1765
rect 3108 1706 4032 1718
rect 3108 1599 3150 1706
rect 3702 1611 4032 1706
rect 4584 1714 5620 1718
rect 4584 1611 5025 1714
rect 5577 1611 5620 1714
rect 3702 1599 5620 1611
rect 3108 1559 5620 1599
rect -24 1444 2488 1499
rect -24 1440 1897 1444
rect -24 1337 18 1440
rect 570 1436 1897 1440
rect 570 1337 908 1436
rect -24 1329 908 1337
rect 1460 1341 1897 1436
rect 2449 1341 2488 1444
rect 1460 1329 2488 1341
rect -24 1297 2488 1329
rect 3108 1452 5620 1507
rect 3108 1448 5029 1452
rect 3108 1345 3150 1448
rect 3702 1444 5029 1448
rect 3702 1345 4040 1444
rect 3108 1337 4040 1345
rect 4592 1349 5029 1444
rect 5581 1349 5620 1452
rect 4592 1337 5620 1349
rect 3108 1305 5620 1337
<< ndiffc >>
rect 7006 1626 7481 1724
rect 7951 1621 8426 1719
rect 8920 1631 9395 1729
rect 7001 1313 7476 1411
rect 7946 1323 8421 1421
rect 8920 1323 9395 1421
rect 1465 167 1689 242
rect 2104 167 2328 242
rect 3168 160 3392 235
rect 3807 160 4031 235
rect 4686 79 4706 99
rect 1469 -117 1693 -24
rect 2085 -117 2309 -24
rect 4757 79 4776 99
rect 3172 -124 3396 -31
rect 3788 -124 4012 -31
<< pdiffc >>
rect 2328 2862 2528 3050
rect 3048 2850 3248 3038
rect 7910 2883 8244 3030
rect 8462 2883 8796 3030
rect 2328 2434 2528 2622
rect 3040 2446 3240 2634
rect 7910 2463 8244 2610
rect 8477 2478 8811 2625
rect 18 1591 570 1698
rect 900 1603 1452 1710
rect 1893 1603 2445 1706
rect 3150 1599 3702 1706
rect 4032 1611 4584 1718
rect 5025 1611 5577 1714
rect 18 1337 570 1440
rect 908 1329 1460 1436
rect 1897 1341 2449 1444
rect 3150 1345 3702 1448
rect 4040 1337 4592 1444
rect 5029 1349 5581 1452
<< psubdiff >>
rect 6942 1215 9464 1254
rect 6942 1117 6996 1215
rect 7471 1117 7951 1215
rect 8426 1117 8925 1215
rect 9400 1117 9464 1215
rect 6942 1078 9464 1117
rect 1394 -222 2396 -195
rect 1394 -338 1457 -222
rect 1685 -225 2396 -222
rect 1685 -338 2085 -225
rect 1394 -341 2085 -338
rect 2313 -341 2396 -225
rect 1394 -397 2396 -341
rect 3097 -229 4099 -202
rect 3097 -345 3160 -229
rect 3388 -232 4099 -229
rect 3388 -345 3788 -232
rect 3097 -348 3788 -345
rect 4016 -348 4099 -232
rect 3097 -398 4099 -348
<< nsubdiff >>
rect 2276 3441 3280 3495
rect 2276 3437 3012 3441
rect 2276 3249 2340 3437
rect 2540 3253 3012 3437
rect 3212 3253 3280 3441
rect 2540 3249 3280 3253
rect 2276 3152 3280 3249
<< psubdiffcont >>
rect 6996 1117 7471 1215
rect 7951 1117 8426 1215
rect 8925 1117 9400 1215
rect 1457 -338 1685 -222
rect 2085 -341 2313 -225
rect 3160 -345 3388 -229
rect 3788 -348 4016 -232
<< nsubdiffcont >>
rect 2340 3249 2540 3437
rect 3012 3253 3212 3441
<< poly >>
rect 5131 2848 5328 2946
rect 5131 2774 5164 2848
rect 3328 2754 5164 2774
rect 2205 2706 2276 2754
rect 3280 2731 5164 2754
rect 5293 2774 5328 2848
rect 5293 2772 7808 2774
rect 5293 2731 7848 2772
rect 3280 2722 7848 2731
rect 8864 2722 8956 2772
rect 3280 2706 7808 2722
rect 3328 2697 7808 2706
rect -417 1630 -170 1662
rect -417 1479 -385 1630
rect -194 1583 -170 1630
rect -194 1551 -75 1583
rect 5782 1662 6029 1670
rect 5782 1599 5830 1662
rect 5678 1559 5830 1599
rect -194 1499 -24 1551
rect 2488 1499 2531 1551
rect 3057 1507 3108 1559
rect 5620 1511 5830 1559
rect 6021 1511 6029 1662
rect 5620 1507 6029 1511
rect -194 1479 -75 1499
rect -417 1463 -75 1479
rect -417 1407 -170 1463
rect 5678 1479 6029 1507
rect 6558 1588 6914 1614
rect 6558 1506 6584 1588
rect 6684 1552 6914 1588
rect 6684 1506 6948 1552
rect 6558 1499 6948 1506
rect 9468 1499 9511 1552
rect 6558 1484 6914 1499
rect 6558 1480 6862 1484
rect 5782 1415 6029 1479
rect 2450 121 3044 144
rect 2450 107 2615 121
rect 1293 51 1401 107
rect 2400 72 2615 107
rect 2664 100 3044 121
rect 2664 72 3104 100
rect 2400 53 3104 72
rect 2400 51 2497 53
rect 2996 44 3104 53
rect 4103 44 4200 100
<< polycont >>
rect 5164 2731 5293 2848
rect -385 1479 -194 1630
rect 5830 1511 6021 1662
rect 6584 1506 6684 1588
rect 2615 72 2664 121
<< ndiffres >>
rect 4676 99 4716 109
rect 4676 79 4686 99
rect 4706 79 4716 99
rect 4676 38 4716 79
rect 4745 99 4786 110
rect 4745 79 4757 99
rect 4776 79 4786 99
rect 4745 70 4786 79
rect 4746 38 4786 70
rect 4676 9 4786 38
<< locali >>
rect 2277 3492 3283 3501
rect 2277 3451 8109 3492
rect 2277 3441 8119 3451
rect 2277 3437 3008 3441
rect 2277 3249 2340 3437
rect 2540 3257 3008 3437
rect 2540 3253 3012 3257
rect 3212 3253 8119 3441
rect 2540 3249 8119 3253
rect 2277 3246 8119 3249
rect 2277 3050 3283 3246
rect 7864 3118 8119 3246
rect 2277 2866 2324 3050
rect 2528 3038 3283 3050
rect 2277 2862 2328 2866
rect 2528 2862 3048 3038
rect 3248 3034 3283 3038
rect 2277 2850 3048 2862
rect 3252 2850 3283 3034
rect 7844 3030 8867 3118
rect 2277 2782 3283 2850
rect 5131 2848 5328 2946
rect 5131 2731 5164 2848
rect 5293 2731 5328 2848
rect 7844 2883 7910 3030
rect 8244 2883 8462 3030
rect 8796 2883 8867 3030
rect 7844 2823 8867 2883
rect 5131 2697 5328 2731
rect 2277 2634 3279 2674
rect 2277 2622 3040 2634
rect 2277 2434 2328 2622
rect 2528 2446 3040 2622
rect 3240 2446 3279 2634
rect 2528 2434 3279 2446
rect 2277 2418 3279 2434
rect 7849 2625 8873 2681
rect 7849 2610 8477 2625
rect 7849 2463 7910 2610
rect 8244 2478 8477 2610
rect 8811 2622 8873 2625
rect 8811 2478 8878 2622
rect 8244 2463 8878 2478
rect 2261 2386 3335 2418
rect 7849 2407 8878 2463
rect 2261 2298 2488 2386
rect 2219 1858 2488 2298
rect 3108 2306 3335 2386
rect 3108 2237 3383 2306
rect 3114 1858 3383 2237
rect 8590 2181 8878 2407
rect 8590 2180 9655 2181
rect 9867 2180 9984 2185
rect 8590 1992 9984 2180
rect 2196 1807 2488 1858
rect 2196 1762 2483 1807
rect -14 1718 2483 1762
rect 3112 1770 3399 1858
rect 3112 1718 5613 1770
rect 8923 1763 9211 1992
rect 9629 1989 9984 1992
rect -14 1710 2481 1718
rect -14 1698 900 1710
rect -425 1630 -154 1662
rect -425 1479 -385 1630
rect -194 1479 -154 1630
rect -14 1591 18 1698
rect 570 1603 900 1698
rect 1452 1706 2481 1710
rect 1452 1603 1893 1706
rect 2445 1603 2481 1706
rect 570 1591 2481 1603
rect -14 1571 2481 1591
rect 3118 1706 4032 1718
rect 3118 1599 3150 1706
rect 3702 1611 4032 1706
rect 4584 1714 5613 1718
rect 4584 1611 5025 1714
rect 5577 1611 5613 1714
rect 6952 1729 9469 1763
rect 6952 1724 8920 1729
rect 3702 1599 5613 1611
rect 3118 1579 5613 1599
rect 5766 1662 6037 1670
rect 5766 1511 5830 1662
rect 6021 1511 6037 1662
rect 6952 1626 7006 1724
rect 7481 1719 8920 1724
rect 7481 1626 7951 1719
rect 6952 1621 7951 1626
rect 8426 1631 8920 1719
rect 9395 1631 9469 1729
rect 8426 1621 9469 1631
rect -425 1407 -154 1479
rect -10 1444 2485 1484
rect -10 1440 1897 1444
rect -10 1337 18 1440
rect 570 1436 1897 1440
rect 570 1337 908 1436
rect -10 1329 908 1337
rect 1460 1341 1897 1436
rect 2449 1341 2485 1444
rect 1460 1329 2485 1341
rect -10 1293 2485 1329
rect 3122 1452 5617 1492
rect 3122 1448 5029 1452
rect 3122 1345 3150 1448
rect 3702 1444 5029 1448
rect 3702 1345 4040 1444
rect 3122 1337 4040 1345
rect 4592 1349 5029 1444
rect 5581 1349 5617 1452
rect 5766 1415 6037 1511
rect 6558 1588 6714 1619
rect 6952 1592 9469 1621
rect 6558 1506 6584 1588
rect 6684 1506 6714 1588
rect 4592 1337 5617 1349
rect 3122 1301 5617 1337
rect 2236 1178 2395 1293
rect 2228 1065 2395 1178
rect 3192 1176 3336 1301
rect 3192 1120 3348 1176
rect 2228 531 2382 1065
rect 3194 781 3348 1120
rect 4670 997 4717 1002
rect 6558 997 6714 1506
rect 6942 1421 9464 1460
rect 6942 1411 7946 1421
rect 6942 1313 7001 1411
rect 7476 1323 7946 1411
rect 8421 1323 8920 1421
rect 9395 1323 9464 1421
rect 7476 1313 9464 1323
rect 6942 1217 9464 1313
rect 6942 1215 7000 1217
rect 7471 1215 9464 1217
rect 6942 1117 6996 1215
rect 7471 1212 7951 1215
rect 7471 1119 7947 1212
rect 7471 1117 7951 1119
rect 8426 1117 8925 1215
rect 9400 1212 9464 1215
rect 9405 1119 9464 1212
rect 9400 1117 9464 1119
rect 6942 1078 9464 1117
rect 4670 924 6718 997
rect 4670 781 4717 924
rect 8618 824 8830 825
rect 9867 824 9984 1989
rect 8618 805 9984 824
rect 7774 792 8238 795
rect 7723 789 8238 792
rect 3194 642 4718 781
rect 6354 775 8238 789
rect 6354 735 7824 775
rect 8176 735 8238 775
rect 8618 765 8643 805
rect 8770 765 9984 805
rect 8618 744 9984 765
rect 8618 738 8850 744
rect 8618 735 8830 738
rect 6354 716 8238 735
rect 2228 459 2717 531
rect 2228 422 2724 459
rect 2228 275 2382 422
rect 1431 253 2382 275
rect 1431 242 2373 253
rect 1431 167 1465 242
rect 1689 167 2104 242
rect 2328 167 2373 242
rect 1431 141 2373 167
rect 2596 121 2724 422
rect 3194 268 3348 642
rect 3134 235 4076 268
rect 3134 160 3168 235
rect 3392 160 3807 235
rect 4031 160 4076 235
rect 3134 134 4076 160
rect 2596 72 2615 121
rect 2664 72 2724 121
rect 4675 99 4717 642
rect 6364 622 6401 716
rect 7723 712 8238 716
rect 7774 710 8238 712
rect 6369 112 6396 622
rect 4792 111 6401 112
rect 4675 89 4686 99
rect 2596 46 2724 72
rect 4676 79 4686 89
rect 4706 89 4717 99
rect 4746 99 6401 111
rect 4706 79 4716 89
rect 4676 69 4716 79
rect 4746 79 4757 99
rect 4776 79 6401 99
rect 4746 76 6401 79
rect 4746 71 4809 76
rect 4746 70 4808 71
rect 7595 39 7692 149
rect 1420 -24 2373 25
rect 1420 -117 1469 -24
rect 1693 -117 2085 -24
rect 2309 -117 2373 -24
rect 1420 -222 2373 -117
rect 1420 -342 1457 -222
rect 1685 -225 2373 -222
rect 1686 -341 2085 -225
rect 2313 -341 2373 -225
rect 1686 -342 2089 -341
rect 2307 -342 2373 -341
rect 1420 -375 2373 -342
rect 3123 -31 4076 18
rect 3123 -124 3172 -31
rect 3396 -124 3788 -31
rect 4012 -124 4076 -31
rect 3123 -229 4076 -124
rect 3123 -345 3160 -229
rect 3388 -232 4076 -229
rect 3393 -342 3785 -232
rect 3388 -345 3788 -342
rect 3123 -348 3788 -345
rect 4016 -348 4076 -232
rect 3123 -382 4076 -348
<< viali >>
rect 2340 3249 2536 3437
rect 3008 3257 3012 3441
rect 3012 3257 3212 3441
rect 2324 2866 2328 3050
rect 2328 2866 2528 3050
rect 3048 2850 3248 3034
rect 3248 2850 3252 3034
rect 7000 1215 7471 1217
rect 7000 1119 7471 1215
rect 7947 1119 7951 1212
rect 7951 1119 8423 1212
rect 8929 1119 9400 1212
rect 9400 1119 9405 1212
rect 7824 735 8176 775
rect 8643 765 8770 805
rect 1457 -338 1685 -225
rect 1685 -338 1686 -225
rect 1457 -342 1686 -338
rect 2089 -341 2307 -225
rect 2089 -342 2307 -341
rect 3164 -342 3388 -232
rect 3388 -342 3393 -232
rect 3785 -342 3788 -232
rect 3788 -342 4014 -232
<< metal1 >>
rect 2237 3441 3311 3485
rect 2237 3437 3008 3441
rect 2237 3249 2340 3437
rect 2536 3257 3008 3437
rect 3212 3257 3311 3441
rect 2536 3249 3311 3257
rect 2237 3050 3311 3249
rect 2237 2866 2324 3050
rect 2528 3034 3311 3050
rect 2528 2866 3048 3034
rect 2237 2850 3048 2866
rect 3252 2850 3311 3034
rect 2237 2810 3311 2850
rect 6908 1239 9498 1450
rect 4356 1217 9498 1239
rect 4356 1119 7000 1217
rect 7471 1212 9498 1217
rect 7471 1119 7947 1212
rect 8423 1119 8929 1212
rect 9405 1119 9498 1212
rect 4356 1097 9498 1119
rect 4356 1057 7009 1097
rect 1340 5 2450 12
rect 1331 -222 4154 5
rect 4364 -222 4477 1057
rect 6802 149 6850 1057
rect 8618 805 8795 828
rect 7782 775 8241 795
rect 7782 735 7824 775
rect 8176 735 8241 775
rect 8618 765 8643 805
rect 8770 765 8795 805
rect 8618 735 8795 765
rect 7782 710 8241 735
rect 6800 146 7548 149
rect 6800 144 7553 146
rect 6800 116 7685 144
rect 6800 62 7620 116
rect 7667 62 7685 116
rect 6800 43 7685 62
rect 6802 19 6850 43
rect 7516 42 7685 43
rect 1331 -225 4477 -222
rect 1331 -342 1457 -225
rect 1686 -342 2089 -225
rect 2307 -232 4477 -225
rect 2307 -342 3164 -232
rect 3393 -342 3785 -232
rect 4014 -342 4477 -232
rect 1331 -366 4477 -342
rect 1340 -372 2450 -366
rect 3044 -377 4477 -366
rect 3044 -379 4154 -377
<< via1 >>
rect 7620 62 7667 116
<< metal2 >>
rect 8765 678 8790 685
rect 7788 675 8242 678
rect 8480 675 8790 678
rect 7693 668 8790 675
rect 7693 667 8788 668
rect 7693 146 8786 667
rect 7593 116 8786 146
rect 7593 62 7620 116
rect 7667 62 8786 116
rect 7593 42 8786 62
rect 7693 -413 8786 42
<< metal3 >>
rect 8620 678 8788 823
rect 8480 675 8790 678
rect 7693 322 8790 675
rect 7693 -413 8786 322
<< mimcap >>
rect 7741 532 8738 632
rect 7741 170 7831 532
rect 8185 170 8738 532
rect 7741 -365 8738 170
<< mimcapcontact >>
rect 7831 170 8185 532
<< metal4 >>
rect 7787 678 8238 793
rect 7787 663 8242 678
rect 7789 532 8242 663
rect 7789 170 7831 532
rect 8185 170 8242 532
rect 7789 107 8242 170
<< labels >>
rlabel locali 2683 61 2702 125 1 vg
rlabel metal1 1715 -359 1771 -221 1 gnd
rlabel locali 3250 439 3300 571 1 vo
rlabel locali -385 1407 -210 1463 1 vinp
rlabel locali 5837 1423 6012 1479 1 vinm
rlabel metal1 2355 3152 2532 3216 1 vdd
rlabel locali 5164 2878 5280 2917 1 vbias
rlabel locali 9876 1436 9970 1481 1 vout
rlabel locali 6713 736 6783 766 1 top
rlabel metal4 7931 716 8004 729 1 top
rlabel metal3 8671 744 8728 759 1 vout
rlabel metal2 7615 126 7660 144 1 gnd
<< end >>
